* C:\Program Files\ADI\LTspice\Draft1.asc
* Input RF Transformer
L1 0 ANT_IN 200µ
L2 0 N004 200µ

* Output RF Transformer
L3 N002 VCC 200µ
L4 0 N001 200µ

* Tuning Capacitor
C1 N004 0 142.32p

* DC Blocking Capacitor
C2 N003 N004 1µ

* RF Tuning Capacitor
C3 VCC N002 142.32p

* DC Biasing Network
R1 VCC N003 47k
R2 N003 0 10k

* Emitter Network
R3 N005 0 220
C4 N005 0 1n

* BC547b Amplifier
Q1 N002 N003 N005 0 BC547B

R_Ant_Res ANT_IN N006 50
R_Mixer N001 0 1k

* Signals & Voltages
B1 N006 0 V=A*(1 + m*sin(2*pi*fm*time)) * sin(2*pi*fc*time)
V1 VCC 0 12

* Models
.model BC547B NPN(IS=2.39E-14 NF=1.008 ISE=3.545E-15 NE=1.541 BF=294.3
+ IKF=0.1357 VAF=63.2 NR=1.004 ISC=6.272E-14 NC=1.243 BR=7.946 IKR=0.1144 
+ VAR=25.9 RB=1 IRB=1.00E-06 RBM=1 RE=0.4683 RC=0.85 XTB=0 EG=1.11 XTI=3 
+ CJE=1.358E-11 VJE=0.65 MJE=0.3279 TF=4.391E-10 XTF=120 VTF=2.643 ITF=0.7495 
+ PTF=0 CJC=3.728E-12 VJC=0.3997 MJC=0.2955 XCJC=0.6193 TR=1.00E-32 CJS=0 
+ VJS=0.75 MJS=0.333 FC=0.9579 Vceo=45 Icrating=100m mfg=NXP)

* Param
.param fc=450k
.param fm=20k
.param m=0.7
.param A=0.1
.tran 1u 1m 0 100n

* Coupling
K1 L1 L2 1
K2 L3 L4 1

.end