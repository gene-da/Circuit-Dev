* Common-Emitter Amplifier Test - Fixed & Verified Version

* Power supply
VCC VCC 0 DC 12

* Input signal (AC only)
Vin VIN 0 AC 1

* Improved bias: sets Vb ~ 2.7V (to allow Ve ≈ 2V for 2mA through 1k)
R1 VCC BIAS 47k
R2 BIAS 0 10k

* DC block and signal injection
CIN VIN BASE 10u

* Transistor
Q1 COLLECTOR BASE EMITTER BC547B

* Collector resistor
RC VCC COLLECTOR 4.7k

* Emitter resistor + bypass cap
RE EMITTER 0 1k
CE EMITTER 0 100u

* Output coupling cap
COUT COLLECTOR OUT 1u

* Output load
RL OUT 0 10k

* BC547B model
.model BC547B NPN(IS=2.39E-14 NF=1.008 ISE=3.545E-15 NE=1.541 BF=294.3 IKF=0.1357 VAF=63.2 NR=1.004 ISC=6.272E-14 NC=1.243 BR=7.946 IKR=0.1144 VAR=25.9 RB=1 IRB=1.00E-06 RBM=1 RE=0.4683 RC=0.85 XTB=0 EG=1.11 XTI=3 CJE=1.358E-11 VJE=0.65 MJE=0.3279 TF=4.391E-10 XTF=120 VTF=2.643 ITF=0.7495 PTF=0 CJC=3.728E-12 VJC=0.3997 MJC=0.2955 XCJC=0.6193 TR=1.00E-32 CJS=0 VJS=0.75 MJS=0.333 FC=0.9579 Vceo=45 Icrating=100m mfg=NXP)

* DC operating point check
.op
.print V(BASE) V(EMITTER) V(COLLECTOR)

* AC sweep (up to 100 MHz is plenty)
.ac dec 100 10 100Meg

.end
